`include "global_params.vh"

module gpr (
    input  clk,
    input  index,
    input  enable,
    output data
);

endmodule
