// general purpose registers
// index
localparam R0 = 8'd0;
localparam R1 = 8'd1;
localparam R2 = 8'd2;
localparam R3 = 8'd3;
localparam R4 = 8'd4;
localparam R5 = 8'd5;
localparam R6 = 8'd6;
localparam R7 = 8'd7;
