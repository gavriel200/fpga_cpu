module alu (
    input  clk,
    output data
);

endmodule
