module interrupt (
    output status
);

endmodule
