module flags (
    input clk
    // input data ?
    // output reg f_carray ??
);

endmodule
