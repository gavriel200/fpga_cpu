module decoder (
    input clk
);

endmodule
